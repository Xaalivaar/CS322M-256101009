module myxor(
    input a,
    input b,
    output y
);

    assign y = a ^ b; // XOR operation
endmodule